//////////////////////////////////////////////////////////////////////
//     design: input_ctrl.v
//////////////////////////////////////////////////////////////////////

// Input controller for each physical input channel: cw/ccw/pe).
// Two single-entry buffers for two virtual channels:(even & odd).
// Accepts on VC that is *external* this cycle:
//     polarity==0 (even cycle): external VC = ODD  -> latch odd, r_out = ~odd_valid
//     polarity==1 (odd  cycle): external VC = EVEN -> latch even, r_out = ~even_valid
// Clear asserted by arbitrator when that VC was forwarded.

`timescale 1ns/1ps

module input_ctrl (
	input  wire        clk,
	input  wire        reset, // active-high synchronous reset
	input  wire        polarity, // indicates if current clk cycle is even (0) or odd (1)

	input  wire        send_in, // send handshaking signal, meaning input valid and should be taken
	output reg         ready_in, // ready handshaking signal, meaning channel is empty and can take data
	input  wire [63:0] data_in, // data input

	// Clear is generated by arbitrator.
	// It is asserted to 1 when arbitrator consumes the data and put into matching output buffer.
	// It is asserted to 0 when arbitrator does not consume the data, i.e. still waiting.
	input  wire        clear_even,
	input  wire        clear_odd,

	// Valid is generated by input_ctrl, meaning the channel is occupied right now.
	// It is asserted to 1 when it accept a packet data.
	// It is asserted to 0 when arbitrator consumes the data via clear.
	output reg         valid_even,
	output reg         valid_odd,

	// Output data for arbitrator.
	output reg  [63:0] data_even,
	output reg  [63:0] data_odd
);

    wire ext_even =  polarity;  // when 1, external is even
    wire ext_odd  = ~polarity;  // when 0, external is odd
    wire can_accept_even = ext_even && !valid_even;
    wire can_accept_odd  = ext_odd  && !valid_odd;

    // This drives me crazy...
    // After several hours of debugging, this seems to be the culprit...
    // ready_in should be driven directly by the current valid_* state, instead of being registered with a non-blocking statement.
    always @(*) begin
        ready_in <= ext_even ? ~valid_even : ~valid_odd;
    end

	always @(posedge clk) begin
		if (reset) begin
			ready_in   <= 1'b1;
			valid_even <= 1'b0;
			valid_odd  <= 1'b0;
			data_even  <= 64'b0;
			data_odd   <= 64'b0;
		end
		else begin
			// If polarity == 1, internal is odd, external is even.
			// If even is not occupied, it is ready for new package.
			// If polarity == 0, internal is even, external is odd.
			// If odd is not occupied, it is ready for new package.
			

			// Latch input if valid and channel empty.
            if (send_in && can_accept_even) begin
                data_even  <= data_in;
                valid_even <= 1'b1;
            end
            if (send_in && can_accept_odd) begin
                data_odd   <= data_in;
                valid_odd  <= 1'b1;
            end

			// If even/odd is consumed in the last cycle: clear == 1'b1,
			// even/odd should no longer be valid
			if (clear_even) valid_even <= 1'b0;
			if (clear_odd)  valid_odd  <= 1'b0;			
		end
	end

endmodule