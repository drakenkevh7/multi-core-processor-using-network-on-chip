//////////////////////////////////////////////////////////////////////
//     design: output_ctrl.v
//////////////////////////////////////////////////////////////////////

// Output controller for each physical output channel: cw/ccw/pe).
// Two single-entry buffers for two virtual channels:(even & odd).
// INTERNAL writes (allocator): only into VC == polarity (even on even, odd on odd).
// EXTERNAL send: VC == ~polarity goes on the wire if valid & r_in.

`timescale 1ns/1ps

module output_ctrl (
	input  wire        clk,
	input  wire        reset, // active-high synchronous reset
	input  wire        polarity, // indicates if current clk cycle is even (0) or odd (1)

	input  wire        ready_out, // ready handshaking signal for output channel.
	output reg         send_out, // send handshaking signal for output channel.
	output reg [63:0] data_out, // data output

	// Data and enable are generated by arbitrator.
	input  wire [63:0] data_even,
	input  wire        en_even,
	input  wire [63:0] data_odd,
	input  wire        en_odd,

	// Let Arbitrator know once data is transmitted.
	output reg         empty_even,
	output reg         empty_odd
);

	// Output buffers 
	reg [63:0] output_buffer_data_even,  output_buffer_data_odd;
    reg        output_buffer_valid_even, output_buffer_valid_odd;

	// Internal even (0) or odd (1)
	// External even (1) or odd (0)
	// Combinational logic for outputs
	always @(*) begin
		data_out = polarity ? output_buffer_data_even : output_buffer_data_odd;
		send_out = polarity ? (output_buffer_valid_even & ready_out) : (output_buffer_valid_odd & ready_out);
		empty_even = !output_buffer_valid_even;
		empty_odd  = !output_buffer_valid_odd;
	end

	always @(posedge clk) begin
		if (reset) begin
			output_buffer_data_even <= 64'b0;
			output_buffer_data_odd  <= 64'b0;
			output_buffer_valid_even <= 1'b0;
			output_buffer_valid_odd  <= 1'b0;
		end
		else begin
			if (polarity) begin
				if (en_odd && !output_buffer_valid_odd) begin
					output_buffer_data_odd <= data_odd;
					output_buffer_valid_odd <= en_odd;
				end
			end
			else begin
				if (en_even && !output_buffer_valid_even) begin
					output_buffer_data_even  <= data_even;
					output_buffer_valid_even <= en_even;
				end
			end

			if (!polarity && output_buffer_data_odd  && ready_out) output_buffer_valid_odd  <= 1'b0;
            if (polarity  && output_buffer_data_even && ready_out) output_buffer_valid_even <= 1'b0;
		end
	end

endmodule